// TCES 330, Spring 2020
// Taras Martynyuk, Ben Mulyarchuk, Kevin Nguyen
// 5/20/2020
// ProjectB
// This is a Verilog description for an 256 x 16 register file

module ControlUnit(reset, clk, data, PC_Out, IR_Out, OutState, NextState, D_Addr, D_Wr,RF_s, RF_W_en, RF_Ra_Addr, RF_Rb_Addr, RF_W_Addr, ALU_s0);
    input logic clk, reset, D_Wr, RF_s, RF_W_en;    // clock, reset, Data write enable, MUX select, Register write enable, ALU select bit  
    output logic [6:0] PC_Out;                              // PC address being sent to Instruction memory
    output logic [15:0] IR_Out, data;                       // Data sent to state machine from Instruction Reg, and data sent into IR from Instruction memory
    output logic [3:0] RF_Ra_Addr, RF_Rb_Addr, RF_W_Addr;   // Addresses for A, B, and write destination within the Register file
    output logic [7:0] D_Addr;                              // address within the Data Memory
    output logic [3:0] OutState, NextState;                 // State of State Machine to be shown on board
    output logic [2:0] ALU_s0;                              // ALU select bit
    logic PC_up, PC_clr, IR_ld;

    //InstMemory (address, clock,	q);
    InstMemory U1(PC_Out, clk, data);

    //StateMachine(reset, data, PC_clr, PC_up, IR_ld, D_addr, D_wr, RF_s, RF_W_addr, RF_W_en, RF_Ra_addr, RF_Rb_addr, CurrentState, NextState);
    StateMachine U2(reset, IR_Out, PC_clr, PC_up, IR_ld, D_addr, D_wr, RF_s, RF_W_addr, RF_W_en, RF_Ra_addr, RF_Rb_addr, OutState, NextState);

    //PC_Counter(clk, up, clear, address);
    PC_Counter U3(clk, PC_up, PC_clr, PC_Out);

    //Instruc_Reg (clk, data, load, out);
    Instruc_Reg U4(clk, data, IR_ld, IR_Out);
endmodule

module ControlUnit_tb();
    logic clk, reset, D_Wr, RF_s, RF_W_en, ALU_s0;   // clock, reset, Data write enable, MUX select, Register write enable, ALU select bit  
    logic [6:0] PC_Out;                              // PC address being sent to Instruction memory
    logic [15:0] IR_Out, data;                       // Data sent to state machine from Instruction Reg, and data sent into IR from Instruction memory
    logic [3:0] RF_Ra_Addr, RF_Rb_Addr, RF_W_Addr;   // Addresses for A, B, and write destination within the Register file
    logic [7:0] D_Addr;                              // address within the Data Memory
    logic [3:0] OutState, NextState;                 // State of State Machine to be shown on board

    ControlUnit DUT(reset, clk, data, PC_Out, IR_Out, OutState, NextState, D_Addr, D_Wr,RF_s, RF_W_en, RF_Ra_Addr, RF_Rb_Addr, RF_W_Addr, ALU_s0);

    always begin        //clock signal
        clk = 0; #10;
        clk = 1; #10;
    end

    initial begin
        reset = 1; #22;
        reset = 0; #22;
        wait (NextState == 1); // NOOP
        $display("Time =%0t PC_Out =%7b Instruction Data =%16b Instruction Register Output =%16b RF_Ra_addr =%4b RF_Rb_Addr =%4b RF_W_Addr =%4b D_Addr =%8b OutState =%4b ALU_s0 =%3b D_Wr =%1b RF_s =%1b RF_W_en =%1b", $time, PC_Out, data, IR_Out, RF_Ra_addr, RF_Rb_Addr, RF_W_Addr, D_Addr, OutState, ALU_s0, D_Wr, RF_s, RF_W_en);
        wait (NextState == 1); // LOAD into data Mem[1] from Reg_File[15]
        $display("Time =%0t PC_Out =%7b Instruction Data =%16b Instruction Register Output =%16b RF_Ra_addr =%4b RF_Rb_Addr =%4b RF_W_Addr =%4b D_Addr =%8b OutState =%4b ALU_s0 =%3b D_Wr =%1b RF_s =%1b RF_W_en =%1b", $time, PC_Out, data, IR_Out, RF_Ra_addr, RF_Rb_Addr, RF_W_Addr, D_Addr, OutState, ALU_s0, D_Wr, RF_s, RF_W_en);        
        wait (NextState == 1); // ADD Reg_File[1] + Reg_File[2] into Reg_File[3]
        $display("Time =%0t PC_Out =%7b Instruction Data =%16b Instruction Register Output =%16b RF_Ra_addr =%4b RF_Rb_Addr =%4b RF_W_Addr =%4b D_Addr =%8b OutState =%4b ALU_s0 =%3b D_Wr =%1b RF_s =%1b RF_W_en =%1b", $time, PC_Out, data, IR_Out, RF_Ra_addr, RF_Rb_Addr, RF_W_Addr, D_Addr, OutState, ALU_s0, D_Wr, RF_s, RF_W_en);
        wait (NextState == 1); // SUB Reg_File[10] - Reg_File[9] into Reg_File[0]
        $display("Time =%0t PC_Out =%7b Instruction Data =%16b Instruction Register Output =%16b RF_Ra_addr =%4b RF_Rb_Addr =%4b RF_W_Addr =%4b D_Addr =%8b OutState =%4b ALU_s0 =%3b D_Wr =%1b RF_s =%1b RF_W_en =%1b", $time, PC_Out, data, IR_Out, RF_Ra_addr, RF_Rb_Addr, RF_W_Addr, D_Addr, OutState, ALU_s0, D_Wr, RF_s, RF_W_en);
        wait (NextState == 1); // STORE Reg_File[4] into data Memory[0]
        $display("Time =%0t PC_Out =%7b Instruction Data =%16b Instruction Register Output =%16b RF_Ra_addr =%4b RF_Rb_Addr =%4b RF_W_Addr =%4b D_Addr =%8b OutState =%4b ALU_s0 =%3b D_Wr =%1b RF_s =%1b RF_W_en =%1b", $time, PC_Out, data, IR_Out, RF_Ra_addr, RF_Rb_Addr, RF_W_Addr, D_Addr, OutState, ALU_s0, D_Wr, RF_s, RF_W_en);
        wait (NextState == 1); // HALT
        $display("Time =%0t PC_Out =%7b Instruction Data =%16b Instruction Register Output =%16b RF_Ra_addr =%4b RF_Rb_Addr =%4b RF_W_Addr =%4b D_Addr =%8b OutState =%4b ALU_s0 =%3b D_Wr =%1b RF_s =%1b RF_W_en =%1b", $time, PC_Out, data, IR_Out, RF_Ra_addr, RF_Rb_Addr, RF_W_Addr, D_Addr, OutState, ALU_s0, D_Wr, RF_s, RF_W_en);
        $stop;
    end
endmodule